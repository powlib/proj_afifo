`timescale 1ns / 1ps

module proj_top();


  //proj_lane #(.W(16),.D(8),.X(3),.ID("LANE0"),.EDBG(0)) l0_inst (
  //  .genclk(),.genrst(),.chkclk(),.chkrst(),.errflg0());

endmodule